
// reset_ff.v - 8-bit resettable D flip-flop

module reset_ff #(parameter WIDTH = 32) (
    input       clk, rst,
    input       [WIDTH-1:0] d,
    output reg  [WIDTH-1:0] q
);

always @(posedge clk or posedge rst) begin
    if (rst) q <= 0;
    else     q <= d;
end

endmodule

